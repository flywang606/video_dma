parameter	DATA_WIDTH	=	32;
parameter	ID_WIDTH	=	3;
parameter	ADDR_WIDTH	=	32;
parameter	LEN_WIDTH	=	8;
parameter	SIZE_WIDTH	=	3;

parameter	BURST_WIDTH	=	2;
parameter	CACHE_WIDTH	=	4;
parameter	PROT_WIDTH	=	3;
parameter	QOS_WIDTH	=	4;
parameter	DATA_WIDTH	=	32;
parameter	ID_WIDTH	=	0;
parameter	RESP_WIDTH	=	2;

//
parameter	LINE_COUNT	 =	16;
parameter	STRIDE_COUNT =	16;

//
parameter	ADDRLSB =	3;//fixed me

parameter 	OUTSTANDING_COUNT = 16;
parameter   MAX_BURST 		  = 3;//fixed me